--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:14:59 11/07/2019
-- Design Name:   
-- Module Name:   E:/xilinx/projects/lab3-4/rs_latch_TB.vhd
-- Project Name:  lab3-4
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: rs_latch
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY rs_latch_TB IS
END rs_latch_TB;
 
ARCHITECTURE behavior OF rs_latch_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT rs_latch
    PORT(
         R : IN  std_logic;
         S : IN  std_logic;
         Q_beh : OUT  std_logic;
         nQ_beh : OUT  std_logic;
         Q_str : OUT  std_logic;
         nQ_str : OUT  std_logic;
         Q_param : OUT  std_logic;
         nQ_param : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal R : std_logic := '0';
   signal S : std_logic := '0';

 	--Outputs
   signal Q_beh : std_logic;
   signal nQ_beh : std_logic;
   signal Q_str : std_logic;
   signal nQ_str : std_logic;
   signal Q_param : std_logic;
   signal nQ_param : std_logic;
	signal ASSERT_SIGNAL: std_logic;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: rs_latch PORT MAP (
          R => R,
          S => S,
          Q_beh => Q_beh,
          nQ_beh => nQ_beh,
          Q_str => Q_str,
          nQ_str => nQ_str,
          Q_param => Q_param,
          nQ_param => nQ_param
        );
		  
	main: process
	begin
	  R <= '0' after 5 ns,    -- s = 1 
	       '1' after 15 ns,   -- s = 0 
			 '0' after 20 ns,   -- s = 0
			 '1' after 25 ns;   -- s = 1
			 
	  S <= '1' after 5 ns,   -- r = 0
	       '0' after 10 ns,  -- r = 0 
			 '1' after 25 ns;  -- r = 1
	  wait;
	end process main;
	
	ASSERT_SIGNAL <= (Q_str xor Q_beh) or (nQ_str xor nQ_beh);
 
END;
